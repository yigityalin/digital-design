`timescale 1ns / 1ps

module two_bit_adder_testbench();
    logic a[1:0], b[1:0], c_in, s[1:0], c_out;
    
    two_bit_adder adder(a, b, c_in, s, c_out);

    initial begin
        a[0] = 0; b[0] = 0; c_in = 0; a[1] = 0; b[1] = 0; #10;
        b[1] = 1;                                         #10;
        a[1] = 1; b[1] = 0;                               #10;
        b[1] = 1;                                         #10;
        c_in = 1; a[1] = 0; b[1] = 0;                     #10;
        b[1] = 1;                                         #10;
        a[1] = 1; b[1] = 0;                               #10;
        b[1] = 1;                                         #10;
        b[0] = 1; c_in = 0; a[1] = 0; b[1] = 0;           #10;
        b[1] = 1;                                         #10;
        a[1] = 1; b[1] = 0;                               #10;
        b[1] = 1;                                         #10;
        c_in = 1; a[1] = 0; b[1] = 0;                     #10;
        b[1] = 1;                                         #10;
        a[1] = 1; b[1] = 0;                               #10;
        b[1] = 1;                                         #10;
        a[0] = 1; b[0] = 0; c_in = 0; a[1] = 0; b[1] = 0; #10;
        b[1] = 1;                                         #10;
        a[1] = 1; b[1] = 0;                               #10;
        b[1] = 1;                                         #10;
        c_in = 1; a[1] = 0; b[1] = 0;                     #10;
        b[1] = 1;                                         #10;
        a[1] = 1; b[1] = 0;                               #10;
        b[1] = 1;                                         #10;
        b[0] = 1; c_in = 0; a[1] = 0; b[1] = 0;           #10;
        b[1] = 1;                                         #10;
        a[1] = 1; b[1] = 0;                               #10;
        b[1] = 1;                                         #10;
        c_in = 1; a[1] = 0; b[1] = 0;                     #10;
        b[1] = 1;                                         #10;
        a[1] = 1; b[1] = 0;                               #10;
        b[1] = 1;                                         #10;
    end
endmodule
